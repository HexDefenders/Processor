module tb_datapath();


endmodule
